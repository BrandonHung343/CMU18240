C:/afs/ece.cmu.edu/class/ee240/bin/RISC240/memory.sv